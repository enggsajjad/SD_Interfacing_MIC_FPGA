library verilog;
use verilog.vl_types.all;
entity spi_interface_tf_v_tf is
end spi_interface_tf_v_tf;
